`timescale 1ns/1ps

// Author : Cernalevschi Cristian
// Project: NN handwritten digit recognition
// File   : The top neural network module (synthesizable)

module top_nn (
    input        clk        ,
    input        reset      ,
    input        enable     ,
    input        oled_ready ,
    input        oled_done  ,
    output       out_valid  ,
    output [3:0] net_data   ,
    output       DONE
);

// Parameters
localparam dataWidth       = 16;
localparam outData         = 10;
localparam outWidth        = $clog2(outData);

// Interconnection wires
wire                   rst_n     ;
wire                   mem_valid ;
wire [dataWidth - 1:0] mem_data  ;
wire                   last      ;
wire                   net_valid ;

// Internal registers
reg  renable        ;
reg  last_done      ;
reg  nn_done        ;
reg  oled_out_valid ;
reg  out_valid_flag ;
reg  oled_done_flag ;

// Assignmets
assign rst_n      = ~reset         ;
assign read_en    = renable        ;
assign out_valid  = oled_out_valid ;
assign DONE       = nn_done        ;

// Enable reading from memory
always @(posedge clk) begin
    if (~rst_n)
        renable <= 1'b0;
    else if (last)
        renable <= 1'b0;
    else if (enable & ~last_done)
        renable <= 1'b1;
end

// Active HIGH - done reading from memory
always @(posedge clk) begin
    if (~rst_n)
        last_done <= 1'b0;
    else if (last)
        last_done <= 1'b1;
end

// Active HIGH - nn generated a result
always @(posedge clk) begin
    if (~rst_n)
        nn_done <= 1'b0;
    else if (renable)
        nn_done <= 1'b0;
    else if (net_valid)
        nn_done <= 1'b1;
end

// Flag that indicates that the result generated by the NN was already be sent in order to be displayed to OLED controller
always @(posedge clk) begin
    if (~rst_n)
        out_valid_flag <= 1'b0;
    else if (nn_done & oled_ready)
        out_valid_flag <= 1'b1;
end

// Generate a write valid pulse to OLED controller when it is ready to receive data and NN also gnerated a result
always @(posedge clk) begin
    if (~rst_n)
        oled_out_valid <= 1'b0;
    else if (nn_done & oled_ready & ~out_valid_flag)
        oled_out_valid <= 1'b1;
    else
        oled_out_valid <= 1'b0;
end

always @(posedge clk) begin
    if (~rst_n)
        oled_done_flag <= 1'b0;
    else if (oled_done)
        oled_done_flag <= 1'b1;
end

// Instantiate the neural network memory
nn_memory #(
    .dataWidth (dataWidth )
) i_nn_memory (
    .clk       (clk       ),
    .rst_n     (rst_n     ),
    .ren       (read_en   ),
    .mem_valid (mem_valid ),
    .mem_data  (mem_data  ),
    .data_last (last      )
);

// Instantiate the neural network core
net #(
    .dataWidth     (dataWidth ),
    .outData       (outData   ),
    .outWidth      (outWidth  )
) i_net (
    .clk           (clk       ),
    .rst_n         (rst_n     ),
    .net_valid     (mem_valid ),
    .net_data      (mem_data  ),
    .net_out_valid (net_valid ),
    .net_out_data  (net_data  )
);
    
endmodule