`timescale 1ns/1ps

// Author : Cernalevschi Cristian
// Project: NN handwritten digit recognition
// File   : Sigmoid activation module

module sigmoid_activation (
    input clk,
    input rst_n,
    input sig_valid,
    input [dataWidth - 1:0] sig_in,
    output [dataWidth - 1:0] sig_out
);

endmodule